module tapped_delay_tdc (
	output [6:0] fine_time,
	input CLK,
    input CAN_logic
);

reg [100:0] Sum = 400'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
wire [100:0] Co /* synthesis keep = 1 */;
reg [100:0] Sum_tmp;
reg [6:0] Sum_num;
reg Ci = 0;
reg Hit;
reg Hit_tmp;

always @(posedge CAN_logic) begin
    Sum_tmp = Sum;
    Hit_tmp = ~Hit;
    if(Sum_tmp[100]==Hit_tmp)Sum_num=100;
    else if(Sum_tmp[99]==Hit_tmp)Sum_num=99;
    else if(Sum_tmp[98]==Hit_tmp)Sum_num=98;
    else if(Sum_tmp[97]==Hit_tmp)Sum_num=97;
    else if(Sum_tmp[96]==Hit_tmp)Sum_num=96;
    else if(Sum_tmp[95]==Hit_tmp)Sum_num=95;
    else if(Sum_tmp[94]==Hit_tmp)Sum_num=94;
    else if(Sum_tmp[93]==Hit_tmp)Sum_num=93;
    else if(Sum_tmp[92]==Hit_tmp)Sum_num=92;
    else if(Sum_tmp[91]==Hit_tmp)Sum_num=91;
    else if(Sum_tmp[90]==Hit_tmp)Sum_num=90;
    else if(Sum_tmp[89]==Hit_tmp)Sum_num=89;
    else if(Sum_tmp[88]==Hit_tmp)Sum_num=88;
    else if(Sum_tmp[87]==Hit_tmp)Sum_num=87;
    else if(Sum_tmp[86]==Hit_tmp)Sum_num=86;
    else if(Sum_tmp[85]==Hit_tmp)Sum_num=85;
    else if(Sum_tmp[84]==Hit_tmp)Sum_num=84;
    else if(Sum_tmp[83]==Hit_tmp)Sum_num=83;
    else if(Sum_tmp[82]==Hit_tmp)Sum_num=82;
    else if(Sum_tmp[81]==Hit_tmp)Sum_num=81;
    else if(Sum_tmp[80]==Hit_tmp)Sum_num=80;
    else if(Sum_tmp[79]==Hit_tmp)Sum_num=79;
    else if(Sum_tmp[78]==Hit_tmp)Sum_num=78;
    else if(Sum_tmp[77]==Hit_tmp)Sum_num=77;
    else if(Sum_tmp[76]==Hit_tmp)Sum_num=76;
    else if(Sum_tmp[75]==Hit_tmp)Sum_num=75;
    else if(Sum_tmp[74]==Hit_tmp)Sum_num=74;
    else if(Sum_tmp[73]==Hit_tmp)Sum_num=73;
    else if(Sum_tmp[72]==Hit_tmp)Sum_num=72;
    else if(Sum_tmp[71]==Hit_tmp)Sum_num=71;
    else if(Sum_tmp[70]==Hit_tmp)Sum_num=70;
    else if(Sum_tmp[69]==Hit_tmp)Sum_num=69;
    else if(Sum_tmp[68]==Hit_tmp)Sum_num=68;
    else if(Sum_tmp[67]==Hit_tmp)Sum_num=67;
    else if(Sum_tmp[66]==Hit_tmp)Sum_num=66;
    else if(Sum_tmp[65]==Hit_tmp)Sum_num=65;
    else if(Sum_tmp[64]==Hit_tmp)Sum_num=64;
    else if(Sum_tmp[63]==Hit_tmp)Sum_num=63;
    else if(Sum_tmp[62]==Hit_tmp)Sum_num=62;
    else if(Sum_tmp[61]==Hit_tmp)Sum_num=61;
    else if(Sum_tmp[60]==Hit_tmp)Sum_num=60;
    else if(Sum_tmp[59]==Hit_tmp)Sum_num=59;
    else if(Sum_tmp[58]==Hit_tmp)Sum_num=58;
    else if(Sum_tmp[57]==Hit_tmp)Sum_num=57;
    else if(Sum_tmp[56]==Hit_tmp)Sum_num=56;
    else if(Sum_tmp[55]==Hit_tmp)Sum_num=55;
    else if(Sum_tmp[54]==Hit_tmp)Sum_num=54;
    else if(Sum_tmp[53]==Hit_tmp)Sum_num=53;
    else if(Sum_tmp[52]==Hit_tmp)Sum_num=52;
    else if(Sum_tmp[51]==Hit_tmp)Sum_num=51;
    else if(Sum_tmp[50]==Hit_tmp)Sum_num=50;
    else if(Sum_tmp[49]==Hit_tmp)Sum_num=49;
    else if(Sum_tmp[48]==Hit_tmp)Sum_num=48;
    else if(Sum_tmp[47]==Hit_tmp)Sum_num=47;
    else if(Sum_tmp[46]==Hit_tmp)Sum_num=46;
    else if(Sum_tmp[45]==Hit_tmp)Sum_num=45;
    else if(Sum_tmp[44]==Hit_tmp)Sum_num=44;
    else if(Sum_tmp[43]==Hit_tmp)Sum_num=43;
    else if(Sum_tmp[42]==Hit_tmp)Sum_num=42;
    else if(Sum_tmp[41]==Hit_tmp)Sum_num=41;
    else if(Sum_tmp[40]==Hit_tmp)Sum_num=40;
    else if(Sum_tmp[39]==Hit_tmp)Sum_num=39;
    else if(Sum_tmp[38]==Hit_tmp)Sum_num=38;
    else if(Sum_tmp[37]==Hit_tmp)Sum_num=37;
    else if(Sum_tmp[36]==Hit_tmp)Sum_num=36;
    else if(Sum_tmp[35]==Hit_tmp)Sum_num=35;
    else if(Sum_tmp[34]==Hit_tmp)Sum_num=34;
    else if(Sum_tmp[33]==Hit_tmp)Sum_num=33;
    else if(Sum_tmp[32]==Hit_tmp)Sum_num=32;
    else if(Sum_tmp[31]==Hit_tmp)Sum_num=31;
    else if(Sum_tmp[30]==Hit_tmp)Sum_num=30;
    else if(Sum_tmp[29]==Hit_tmp)Sum_num=29;
    else if(Sum_tmp[28]==Hit_tmp)Sum_num=28;
    else if(Sum_tmp[27]==Hit_tmp)Sum_num=27;
    else if(Sum_tmp[26]==Hit_tmp)Sum_num=26;
    else if(Sum_tmp[25]==Hit_tmp)Sum_num=25;
    else if(Sum_tmp[24]==Hit_tmp)Sum_num=24;
    else if(Sum_tmp[23]==Hit_tmp)Sum_num=23;
    else if(Sum_tmp[22]==Hit_tmp)Sum_num=22;
    else if(Sum_tmp[21]==Hit_tmp)Sum_num=21;
    else if(Sum_tmp[20]==Hit_tmp)Sum_num=20;
    else if(Sum_tmp[19]==Hit_tmp)Sum_num=19;
    else if(Sum_tmp[18]==Hit_tmp)Sum_num=18;
    else if(Sum_tmp[17]==Hit_tmp)Sum_num=17;
    else if(Sum_tmp[16]==Hit_tmp)Sum_num=16;
    else if(Sum_tmp[15]==Hit_tmp)Sum_num=15;
    else if(Sum_tmp[14]==Hit_tmp)Sum_num=14;
    else if(Sum_tmp[13]==Hit_tmp)Sum_num=13;
    else if(Sum_tmp[12]==Hit_tmp)Sum_num=12;
    else if(Sum_tmp[11]==Hit_tmp)Sum_num=11;
    else if(Sum_tmp[10]==Hit_tmp)Sum_num=10;
    else if(Sum_tmp[9]==Hit_tmp)Sum_num=9;
    else if(Sum_tmp[8]==Hit_tmp)Sum_num=8;
    else if(Sum_tmp[7]==Hit_tmp)Sum_num=7;
    else if(Sum_tmp[6]==Hit_tmp)Sum_num=6;
    else if(Sum_tmp[5]==Hit_tmp)Sum_num=5;
    else if(Sum_tmp[4]==Hit_tmp)Sum_num=4;
    else if(Sum_tmp[3]==Hit_tmp)Sum_num=3;
    else if(Sum_tmp[2]==Hit_tmp)Sum_num=2;
    else if(Sum_tmp[1]==Hit_tmp)Sum_num=1;
    else Sum_num=0;
end

adder adder_0(.Sum(Sum[0]), .Co(Co[0]), .A(1), .B(Hit), .Ci(Ci));
adder adder_1(.Sum(Sum[1]), .Co(Co[1]), .A(1), .B(0), .Ci(Co[0]));
adder adder_2(.Sum(Sum[2]), .Co(Co[2]), .A(1), .B(0), .Ci(Co[1]));
adder adder_3(.Sum(Sum[3]), .Co(Co[3]), .A(1), .B(0), .Ci(Co[2]));
adder adder_4(.Sum(Sum[4]), .Co(Co[4]), .A(1), .B(0), .Ci(Co[3]));
adder adder_5(.Sum(Sum[5]), .Co(Co[5]), .A(1), .B(0), .Ci(Co[4]));
adder adder_6(.Sum(Sum[6]), .Co(Co[6]), .A(1), .B(0), .Ci(Co[5]));
adder adder_7(.Sum(Sum[7]), .Co(Co[7]), .A(1), .B(0), .Ci(Co[6]));
adder adder_8(.Sum(Sum[8]), .Co(Co[8]), .A(1), .B(0), .Ci(Co[7]));
adder adder_9(.Sum(Sum[9]), .Co(Co[9]), .A(1), .B(0), .Ci(Co[8]));
adder adder_10(.Sum(Sum[10]), .Co(Co[10]), .A(1), .B(0), .Ci(Co[9]));
adder adder_11(.Sum(Sum[11]), .Co(Co[11]), .A(1), .B(0), .Ci(Co[10]));
adder adder_12(.Sum(Sum[12]), .Co(Co[12]), .A(1), .B(0), .Ci(Co[11]));
adder adder_13(.Sum(Sum[13]), .Co(Co[13]), .A(1), .B(0), .Ci(Co[12]));
adder adder_14(.Sum(Sum[14]), .Co(Co[14]), .A(1), .B(0), .Ci(Co[13]));
adder adder_15(.Sum(Sum[15]), .Co(Co[15]), .A(1), .B(0), .Ci(Co[14]));
adder adder_16(.Sum(Sum[16]), .Co(Co[16]), .A(1), .B(0), .Ci(Co[15]));
adder adder_17(.Sum(Sum[17]), .Co(Co[17]), .A(1), .B(0), .Ci(Co[16]));
adder adder_18(.Sum(Sum[18]), .Co(Co[18]), .A(1), .B(0), .Ci(Co[17]));
adder adder_19(.Sum(Sum[19]), .Co(Co[19]), .A(1), .B(0), .Ci(Co[18]));
adder adder_20(.Sum(Sum[20]), .Co(Co[20]), .A(1), .B(0), .Ci(Co[19]));
adder adder_21(.Sum(Sum[21]), .Co(Co[21]), .A(1), .B(0), .Ci(Co[20]));
adder adder_22(.Sum(Sum[22]), .Co(Co[22]), .A(1), .B(0), .Ci(Co[21]));
adder adder_23(.Sum(Sum[23]), .Co(Co[23]), .A(1), .B(0), .Ci(Co[22]));
adder adder_24(.Sum(Sum[24]), .Co(Co[24]), .A(1), .B(0), .Ci(Co[23]));
adder adder_25(.Sum(Sum[25]), .Co(Co[25]), .A(1), .B(0), .Ci(Co[24]));
adder adder_26(.Sum(Sum[26]), .Co(Co[26]), .A(1), .B(0), .Ci(Co[25]));
adder adder_27(.Sum(Sum[27]), .Co(Co[27]), .A(1), .B(0), .Ci(Co[26]));
adder adder_28(.Sum(Sum[28]), .Co(Co[28]), .A(1), .B(0), .Ci(Co[27]));
adder adder_29(.Sum(Sum[29]), .Co(Co[29]), .A(1), .B(0), .Ci(Co[28]));
adder adder_30(.Sum(Sum[30]), .Co(Co[30]), .A(1), .B(0), .Ci(Co[29]));
adder adder_31(.Sum(Sum[31]), .Co(Co[31]), .A(1), .B(0), .Ci(Co[30]));
adder adder_32(.Sum(Sum[32]), .Co(Co[32]), .A(1), .B(0), .Ci(Co[31]));
adder adder_33(.Sum(Sum[33]), .Co(Co[33]), .A(1), .B(0), .Ci(Co[32]));
adder adder_34(.Sum(Sum[34]), .Co(Co[34]), .A(1), .B(0), .Ci(Co[33]));
adder adder_35(.Sum(Sum[35]), .Co(Co[35]), .A(1), .B(0), .Ci(Co[34]));
adder adder_36(.Sum(Sum[36]), .Co(Co[36]), .A(1), .B(0), .Ci(Co[35]));
adder adder_37(.Sum(Sum[37]), .Co(Co[37]), .A(1), .B(0), .Ci(Co[36]));
adder adder_38(.Sum(Sum[38]), .Co(Co[38]), .A(1), .B(0), .Ci(Co[37]));
adder adder_39(.Sum(Sum[39]), .Co(Co[39]), .A(1), .B(0), .Ci(Co[38]));
adder adder_40(.Sum(Sum[40]), .Co(Co[40]), .A(1), .B(0), .Ci(Co[39]));
adder adder_41(.Sum(Sum[41]), .Co(Co[41]), .A(1), .B(0), .Ci(Co[40]));
adder adder_42(.Sum(Sum[42]), .Co(Co[42]), .A(1), .B(0), .Ci(Co[41]));
adder adder_43(.Sum(Sum[43]), .Co(Co[43]), .A(1), .B(0), .Ci(Co[42]));
adder adder_44(.Sum(Sum[44]), .Co(Co[44]), .A(1), .B(0), .Ci(Co[43]));
adder adder_45(.Sum(Sum[45]), .Co(Co[45]), .A(1), .B(0), .Ci(Co[44]));
adder adder_46(.Sum(Sum[46]), .Co(Co[46]), .A(1), .B(0), .Ci(Co[45]));
adder adder_47(.Sum(Sum[47]), .Co(Co[47]), .A(1), .B(0), .Ci(Co[46]));
adder adder_48(.Sum(Sum[48]), .Co(Co[48]), .A(1), .B(0), .Ci(Co[47]));
adder adder_49(.Sum(Sum[49]), .Co(Co[49]), .A(1), .B(0), .Ci(Co[48]));
adder adder_50(.Sum(Sum[50]), .Co(Co[50]), .A(1), .B(0), .Ci(Co[49]));
adder adder_51(.Sum(Sum[51]), .Co(Co[51]), .A(1), .B(0), .Ci(Co[50]));
adder adder_52(.Sum(Sum[52]), .Co(Co[52]), .A(1), .B(0), .Ci(Co[51]));
adder adder_53(.Sum(Sum[53]), .Co(Co[53]), .A(1), .B(0), .Ci(Co[52]));
adder adder_54(.Sum(Sum[54]), .Co(Co[54]), .A(1), .B(0), .Ci(Co[53]));
adder adder_55(.Sum(Sum[55]), .Co(Co[55]), .A(1), .B(0), .Ci(Co[54]));
adder adder_56(.Sum(Sum[56]), .Co(Co[56]), .A(1), .B(0), .Ci(Co[55]));
adder adder_57(.Sum(Sum[57]), .Co(Co[57]), .A(1), .B(0), .Ci(Co[56]));
adder adder_58(.Sum(Sum[58]), .Co(Co[58]), .A(1), .B(0), .Ci(Co[57]));
adder adder_59(.Sum(Sum[59]), .Co(Co[59]), .A(1), .B(0), .Ci(Co[58]));
adder adder_60(.Sum(Sum[60]), .Co(Co[60]), .A(1), .B(0), .Ci(Co[59]));
adder adder_61(.Sum(Sum[61]), .Co(Co[61]), .A(1), .B(0), .Ci(Co[60]));
adder adder_62(.Sum(Sum[62]), .Co(Co[62]), .A(1), .B(0), .Ci(Co[61]));
adder adder_63(.Sum(Sum[63]), .Co(Co[63]), .A(1), .B(0), .Ci(Co[62]));
adder adder_64(.Sum(Sum[64]), .Co(Co[64]), .A(1), .B(0), .Ci(Co[63]));
adder adder_65(.Sum(Sum[65]), .Co(Co[65]), .A(1), .B(0), .Ci(Co[64]));
adder adder_66(.Sum(Sum[66]), .Co(Co[66]), .A(1), .B(0), .Ci(Co[65]));
adder adder_67(.Sum(Sum[67]), .Co(Co[67]), .A(1), .B(0), .Ci(Co[66]));
adder adder_68(.Sum(Sum[68]), .Co(Co[68]), .A(1), .B(0), .Ci(Co[67]));
adder adder_69(.Sum(Sum[69]), .Co(Co[69]), .A(1), .B(0), .Ci(Co[68]));
adder adder_70(.Sum(Sum[70]), .Co(Co[70]), .A(1), .B(0), .Ci(Co[69]));
adder adder_71(.Sum(Sum[71]), .Co(Co[71]), .A(1), .B(0), .Ci(Co[70]));
adder adder_72(.Sum(Sum[72]), .Co(Co[72]), .A(1), .B(0), .Ci(Co[71]));
adder adder_73(.Sum(Sum[73]), .Co(Co[73]), .A(1), .B(0), .Ci(Co[72]));
adder adder_74(.Sum(Sum[74]), .Co(Co[74]), .A(1), .B(0), .Ci(Co[73]));
adder adder_75(.Sum(Sum[75]), .Co(Co[75]), .A(1), .B(0), .Ci(Co[74]));
adder adder_76(.Sum(Sum[76]), .Co(Co[76]), .A(1), .B(0), .Ci(Co[75]));
adder adder_77(.Sum(Sum[77]), .Co(Co[77]), .A(1), .B(0), .Ci(Co[76]));
adder adder_78(.Sum(Sum[78]), .Co(Co[78]), .A(1), .B(0), .Ci(Co[77]));
adder adder_79(.Sum(Sum[79]), .Co(Co[79]), .A(1), .B(0), .Ci(Co[78]));
adder adder_80(.Sum(Sum[80]), .Co(Co[80]), .A(1), .B(0), .Ci(Co[79]));
adder adder_81(.Sum(Sum[81]), .Co(Co[81]), .A(1), .B(0), .Ci(Co[80]));
adder adder_82(.Sum(Sum[82]), .Co(Co[82]), .A(1), .B(0), .Ci(Co[81]));
adder adder_83(.Sum(Sum[83]), .Co(Co[83]), .A(1), .B(0), .Ci(Co[82]));
adder adder_84(.Sum(Sum[84]), .Co(Co[84]), .A(1), .B(0), .Ci(Co[83]));
adder adder_85(.Sum(Sum[85]), .Co(Co[85]), .A(1), .B(0), .Ci(Co[84]));
adder adder_86(.Sum(Sum[86]), .Co(Co[86]), .A(1), .B(0), .Ci(Co[85]));
adder adder_87(.Sum(Sum[87]), .Co(Co[87]), .A(1), .B(0), .Ci(Co[86]));
adder adder_88(.Sum(Sum[88]), .Co(Co[88]), .A(1), .B(0), .Ci(Co[87]));
adder adder_89(.Sum(Sum[89]), .Co(Co[89]), .A(1), .B(0), .Ci(Co[88]));
adder adder_90(.Sum(Sum[90]), .Co(Co[90]), .A(1), .B(0), .Ci(Co[89]));
adder adder_91(.Sum(Sum[91]), .Co(Co[91]), .A(1), .B(0), .Ci(Co[90]));
adder adder_92(.Sum(Sum[92]), .Co(Co[92]), .A(1), .B(0), .Ci(Co[91]));
adder adder_93(.Sum(Sum[93]), .Co(Co[93]), .A(1), .B(0), .Ci(Co[92]));
adder adder_94(.Sum(Sum[94]), .Co(Co[94]), .A(1), .B(0), .Ci(Co[93]));
adder adder_95(.Sum(Sum[95]), .Co(Co[95]), .A(1), .B(0), .Ci(Co[94]));
adder adder_96(.Sum(Sum[96]), .Co(Co[96]), .A(1), .B(0), .Ci(Co[95]));
adder adder_97(.Sum(Sum[97]), .Co(Co[97]), .A(1), .B(0), .Ci(Co[96]));
adder adder_98(.Sum(Sum[98]), .Co(Co[98]), .A(1), .B(0), .Ci(Co[97]));
adder adder_99(.Sum(Sum[99]), .Co(Co[99]), .A(1), .B(0), .Ci(Co[98]));
adder adder_100(.Sum(Sum[100]), .Co(Co[100]), .A(1), .B(0), .Ci(Co[99]));

always @(posedge CLK) begin
    if (Hit==0) Hit <= 1;
    else Hit <= 0;
end

assign fine_time[6:0] = Sum_num[6:0];

endmodule

